library ieee;
use     ieee.std_logic_1164.all;

entity audio_dsp_top is
port (
);
end audio_dsp_top;

architecture rtl of audio_dsp_top is

begin

end rtl;
